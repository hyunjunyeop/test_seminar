module sadfsadf (
    ports
);
    
endmodule


always @( * )) begin
    
end

always @(dddd) begin
    
end